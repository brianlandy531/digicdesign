* Example circuit file for simulating PEX

.OPTION DOTNODE
.HIER /


.INCLUDE "/home/bxl1703/Pyxis_SPT_HEP/ic_projects/Pyxis_SPT/digicdesign/miniALU/miniALU.cal/miniALU.pex.netlist"

.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_33
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_lwt
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_hwt
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_BIP
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_BIP_NPN
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo DIO
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo DIO_33
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_RES
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo MOS_CAP
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/res.spi res_t


* - Instantiate your parasitic netlist and add the load capacitor
** FORMAT : 
* XLAYOUT [all inputs as listed by the ".subckt" line in the included netlist, in the order that they appear there] [name of the subcircuit as listed in the included netlist]
XLAYOUT COUT OUTPUT[0] INPUT1[0] CONTROL[0] CONTROL[1] INPUT2[0] MINIALU

**--GROUND


**--COUT S0 0 120f
**--COUT S1 0 120f
**--COUT S2 0 120f
**--COUT S3 0 120f
**--COUT COUT 0 120f

**--COUT S0 0 120f
**--COUT S1 0 120f
**--COUT S2 0 120f
**--COUT S3 0 120f


COUT COUT 0 120f

COUT OUTPUT[0] 0 120f



* - Analysis Setup - DC sweep
* FORMAT : .DC [name] [low] [high] [step]
* .DC VFORCE__VIN 0 1.08 0.01

* - Analysis Setup - Trans
* FORMAT : .TRAN [start time] [end time] [time step]
** .TRAN 0 10000n 0.001n
.TRAN 0 10000n 0.001n


* --- Forces
* FORMAT -- PULSE : [name] [port] [reference (0 means ground)] PULSE [low] [high] [delay] [fall time] [rise time] [pulse width] [period]
*
* FORMAT -- DC    : [name] [port] [reference (0 means ground)] DC [voltage]
*
** VFORCE__Vin VIN 0 PULSE (0 1.08 100n 0.1n 0.1n 50n 200n)


**--VFORCE__B0 B0 0 pattern 1.08 0 50n .01n .01n 100n 011 R
**--VFORCE__B1 B1 0 pattern 1.08 0 50n .01n .01n 100n 010 R
**--VFORCE__B2 B2 0 pattern 1.08 0 50n .01n .01n 100n 011 R
**--VFORCE__B3 B3 0 pattern 1.08 0 50n .01n .01n 100n 000 R


**--VFORCE__A0 A0 0 pattern 1.08 0 50n .01n .01n 100n 111 R
**--VFORCE__A1 A1 0 pattern 1.08 0 50n .01n .01n 100n 110 R
**--VFORCE__A2 A2 0 pattern 1.08 0 50n .01n .01n 100n 101 R
**--VFORCE__A3 A3 0 pattern 1.08 0 50n .01n .01n 100n 110 R


**--VFORCE__B0 B0 0 pattern 1.08 0 50n .01n .01n 100n 011 R
**--VFORCE__B1 B1 0 pattern 1.08 0 50n .01n .01n 100n 010 R
**--VFORCE__B2 B2 0 pattern 1.08 0 50n .01n .01n 100n 011 R
**--VFORCE__B3 B3 0 pattern 1.08 0 50n .01n .01n 100n 000 R


VFORCE__VDD VDD 0 DC 1.08
VFORCE__VSS VSS 0 DC 0


** control 00 to 01 to 10 to 11

**00 and 
**01 or 
**10 add 
**11 sub

** each test case will have a zero out period in between
** zero out
** control_0 - 0
** control_1 - 0
** Input2_0 - 0
** Input1_0 - 0




VFORCE__CONTROL[1] CONTROL[1] 0 pattern 1.08 0 50n .01n .01n 100n 0011111111 R
VFORCE__CONTROL[0] CONTROL[0] 0 pattern 1.08 0 50n .01n .01n 100n 0100001111 R

VFORCE__INPUT1[0] INPUT1[0] 0 pattern 1.08 0 50n .01n .01n 100n   1101010101 R
VFORCE__INPUT2[0] INPUT2[0] 0 pattern 1.08 0 50n .01n .01n 100n   0000110011 R

.measure tran static_pwr_hi AVG power from=144.629ns to=248.888ns
.measure tran static_pwr_low AVG power from=283.050ns to=346.610ns

.measure tran inst_pwr MAX power from=0ns to=10000ns

* --- Waveform Outputs
*.PLOT DC V(VIN)
*.PLOT DC V(VOUT)

.PLOT TRAN V(CONTROL[0])
.PLOT TRAN V(CONTROL[1])


.PLOT TRAN V(INPUT1[0])
.PLOT TRAN V(INPUT2[0])
.PLOT TRAN V(OUTPUT[0])

.PLOT TRAN V(COUT)

* --- Params
.TEMP 125


