* SPICE NETLIST
***************************************

.SUBCKT mimcap_g13 plus minus
.ENDS
***************************************
.SUBCKT spiral_inductor_lvs pos neg
.ENDS
***************************************
.SUBCKT mirroradder Vdd GROUND S Cout B Cin A
** N=75 EP=7 IP=0 FDC=28
* PORT Vdd Vdd -1083070 648225 metal1
* PORT GROUND GROUND -1082458 637420 metal1
* PORT S S -1049253 642377 metal1
* PORT Cout Cout -1049368 643362 metal1
* PORT B B -1080430 643400 metal1
* PORT Cin Cin -1078015 643390 metal1
* PORT A A -1082915 643390 metal1
M0 GROUND A 8 GROUND nmos L=1.3e-07 W=5.2e-07 $X=-1082140 $Y=640015 $D=19
M1 8 B GROUND GROUND nmos L=1.3e-07 W=5.2e-07 $X=-1079680 $Y=640015 $D=19
M2 9 Cin 8 GROUND nmos L=1.3e-07 W=5.2e-07 $X=-1077230 $Y=640015 $D=19
M3 10 A 9 GROUND nmos L=1.3e-07 W=5.2e-07 $X=-1074800 $Y=640015 $D=19
M4 GROUND B 10 GROUND nmos L=1.3e-07 W=5.2e-07 $X=-1072320 $Y=640015 $D=19
M5 11 Cin GROUND GROUND nmos L=1.3e-07 W=6.5e-07 $X=-1069890 $Y=639945 $D=19
M6 GROUND B 11 GROUND nmos L=1.3e-07 W=6.5e-07 $X=-1067440 $Y=639945 $D=19
M7 11 A GROUND GROUND nmos L=1.3e-07 W=6.5e-07 $X=-1064990 $Y=639945 $D=19
M8 12 9 11 GROUND nmos L=1.3e-07 W=6.5e-07 $X=-1062545 $Y=639945 $D=19
M9 13 Cin 12 GROUND nmos L=1.3e-07 W=7e-07 $X=-1060090 $Y=639895 $D=19
M10 14 B 13 GROUND nmos L=1.3e-07 W=7e-07 $X=-1057640 $Y=639895 $D=19
M11 GROUND A 14 GROUND nmos L=1.3e-07 W=7e-07 $X=-1055190 $Y=639895 $D=19
M12 S 12 GROUND GROUND nmos L=1.3e-07 W=2.6e-07 $X=-1052740 $Y=640335 $D=19
M13 Cout 9 GROUND GROUND nmos L=1.3e-07 W=2.6e-07 $X=-1050290 $Y=640335 $D=19
M14 Vdd A 15 Vdd pmos L=1.3e-07 W=1.04e-06 $X=-1082140 $Y=644635 $D=25
M15 15 B Vdd Vdd pmos L=1.3e-07 W=1.04e-06 $X=-1079680 $Y=644635 $D=25
M16 9 Cin 15 Vdd pmos L=1.3e-07 W=1.04e-06 $X=-1077230 $Y=644635 $D=25
M17 25 A 9 Vdd pmos L=1.3e-07 W=1.04e-06 $X=-1074800 $Y=644635 $D=25
M18 Vdd B 25 Vdd pmos L=1.3e-07 W=1.04e-06 $X=-1072320 $Y=644635 $D=25
M19 29 Cin Vdd Vdd pmos L=1.3e-07 W=1.3e-06 $X=-1069890 $Y=644695 $D=25
M20 Vdd B 29 Vdd pmos L=1.3e-07 W=1.3e-06 $X=-1067440 $Y=644695 $D=25
M21 29 A Vdd Vdd pmos L=1.3e-07 W=1.3e-06 $X=-1064990 $Y=644695 $D=25
M22 12 9 29 Vdd pmos L=1.3e-07 W=1.3e-06 $X=-1062545 $Y=644695 $D=25
M23 38 Cin 12 Vdd pmos L=1.3e-07 W=1.56e-06 $X=-1060090 $Y=644695 $D=25
M24 41 B 38 Vdd pmos L=1.3e-07 W=1.56e-06 $X=-1057640 $Y=644695 $D=25
M25 Vdd A 41 Vdd pmos L=1.3e-07 W=1.56e-06 $X=-1055190 $Y=644695 $D=25
M26 S 12 Vdd Vdd pmos L=1.3e-07 W=5.2e-07 $X=-1052740 $Y=644695 $D=25
M27 Cout 9 Vdd Vdd pmos L=1.3e-07 W=5.2e-07 $X=-1050290 $Y=644695 $D=25
.ENDS
***************************************
.SUBCKT 4bitripplecarry B0 Cin0 A0 S0 A1 B1 S1 B2 A2 S2 B3 A3 VDD GROUND Cout S3
** N=19 EP=16 IP=28 FDC=112
* PORT B0 B0 -2187988 1305752 metal1
* PORT Cin0 Cin0 -2188015 1304985 metal1
* PORT A0 A0 -2187930 1306822 metal1
* PORT S0 S0 -2152895 1305572 metal1
* PORT A1 A1 -2145313 1306855 metal1
* PORT B1 B1 -2145315 1305727 metal1
* PORT S1 S1 -2110403 1305645 metal1
* PORT B2 B2 -2106385 1305672 metal1
* PORT A2 A2 -2106328 1306762 metal1
* PORT S2 S2 -2071590 1305495 metal1
* PORT B3 B3 -2068900 1305845 metal1
* PORT A3 A3 -2068640 1306795 metal1
* PORT VDD VDD -2187370 1313947 metal1
* PORT GROUND GROUND -2185188 1299397 metal1
* PORT Cout Cout -2034030 1306627 metal1
* PORT S3 S3 -2033920 1305542 metal1
X0 VDD GROUND S0 6 B0 Cin0 A0 mirroradder $T=-1104290 663250 0 0 $X=-2188065 $Y=1300080
X1 VDD GROUND S1 9 B1 6 A1 mirroradder $T=-1061620 663250 0 0 $X=-2145395 $Y=1300080
X2 VDD GROUND S2 13 B2 9 A2 mirroradder $T=-1022755 663150 0 0 $X=-2106530 $Y=1299980
X3 VDD GROUND S3 Cout B3 13 A3 mirroradder $T=-985255 663225 0 0 $X=-2069030 $Y=1300055
.ENDS
***************************************
