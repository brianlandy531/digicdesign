* SPICE NETLIST
***************************************

.SUBCKT mimcap_g13 plus minus
.ENDS
***************************************
.SUBCKT spiral_inductor_lvs pos neg
.ENDS
***************************************
.SUBCKT inv01 VSS VDD Y A
** N=4 EP=4 IP=0 FDC=2
* PORT VSS VSS 980 350 metal1
* PORT VDD VDD 980 8050 metal1
* PORT Y Y 1435 3675 metal1
* PORT A A 805 3675 metal1
M0 Y A VSS VSS nmos L=1.4e-07 W=3.5e-07 $X=910 $Y=1820 $D=19
M1 Y A VDD VDD pmos L=1.4e-07 W=7.7e-07 $X=910 $Y=5600 $D=25
.ENDS
***************************************
.SUBCKT aoi222 VDD Y 3 A0 A1 B1 B0 C0 C1
** N=14 EP=9 IP=0 FDC=12
* PORT VDD VDD 2695 8050 metal1
* PORT Y Y 4375 3675 metal1
* PORT A0 A0 560 3675 metal1
* PORT A1 A1 1190 3045 metal1
* PORT B1 B1 1820 4305 metal1
* PORT B0 B0 2450 3675 metal1
* PORT C0 C0 3080 3045 metal1
* PORT C1 C1 3745 4305 metal1
M0 10 A0 Y 3 nmos L=1.4e-07 W=9.1e-07 $X=770 $Y=1190 $D=19
M1 3 A1 10 3 nmos L=1.4e-07 W=9.1e-07 $X=1190 $Y=1190 $D=19
M2 11 B1 3 3 nmos L=1.4e-07 W=7.7e-07 $X=1785 $Y=1330 $D=19
M3 Y B0 11 3 nmos L=1.4e-07 W=7.7e-07 $X=2205 $Y=1330 $D=19
M4 12 C0 Y 3 nmos L=1.4e-07 W=7.7e-07 $X=2765 $Y=1330 $D=19
M5 3 C1 12 3 nmos L=1.4e-07 W=7.7e-07 $X=3185 $Y=1330 $D=19
M6 VDD A0 13 VDD pmos L=1.4e-07 W=1.82e-06 $X=770 $Y=5390 $D=25
M7 13 A1 VDD VDD pmos L=1.4e-07 W=1.82e-06 $X=1330 $Y=5390 $D=25
M8 14 B1 13 VDD pmos L=1.4e-07 W=1.61e-06 $X=1925 $Y=5390 $D=25
M9 13 B0 14 VDD pmos L=1.4e-07 W=1.61e-06 $X=2485 $Y=5390 $D=25
M10 Y C0 14 VDD pmos L=1.4e-07 W=1.61e-06 $X=3605 $Y=5390 $D=25
M11 14 C1 Y VDD pmos L=1.4e-07 W=1.61e-06 $X=4165 $Y=5390 $D=25
.ENDS
***************************************
.SUBCKT nand02 VSS Y VDD A1 A0
** N=6 EP=5 IP=0 FDC=4
* PORT VSS VSS 1225 350 metal1
* PORT Y Y 1925 3675 metal1
* PORT VDD VDD 1225 8050 metal1
* PORT A1 A1 665 3675 metal1
* PORT A0 A0 1295 4305 metal1
M0 6 A1 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=875 $Y=1190 $D=19
M1 Y A0 6 VSS nmos L=1.4e-07 W=7.7e-07 $X=1295 $Y=1190 $D=19
M2 Y A1 VDD VDD pmos L=1.4e-07 W=1.05e-06 $X=875 $Y=6160 $D=25
M3 VDD A0 Y VDD pmos L=1.4e-07 W=1.05e-06 $X=1435 $Y=6160 $D=25
.ENDS
***************************************
.SUBCKT aoi21 VSS VDD Y A1 A0 B0
** N=8 EP=6 IP=0 FDC=6
* PORT VSS VSS 1470 350 metal1
* PORT VDD VDD 1470 8050 metal1
* PORT Y Y 2485 3675 metal1
* PORT A1 A1 560 3675 metal1
* PORT A0 A0 1190 3045 metal1
* PORT B0 B0 1855 4305 metal1
M0 7 A1 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=805 $Y=1170 $D=19
M1 Y A0 7 VSS nmos L=1.4e-07 W=7.7e-07 $X=1225 $Y=1170 $D=19
M2 VSS B0 Y VSS nmos L=1.4e-07 W=3.5e-07 $X=1820 $Y=1590 $D=19
M3 VDD A1 8 VDD pmos L=1.4e-07 W=1.19e-06 $X=805 $Y=6020 $D=25
M4 8 A0 VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=1365 $Y=6020 $D=25
M5 Y B0 8 VDD pmos L=1.4e-07 W=1.19e-06 $X=1925 $Y=6020 $D=25
.ENDS
***************************************
.SUBCKT xnor2 VDD VSS Y A0 A1
** N=9 EP=5 IP=0 FDC=10
* PORT VDD VDD 2450 8050 metal1
* PORT VSS VSS 2450 350 metal1
* PORT Y Y 3955 3675 metal1
* PORT A0 A0 980 3675 metal1
* PORT A1 A1 2555 3675 metal1
M0 7 A0 6 VSS nmos L=1.4e-07 W=7.7e-07 $X=805 $Y=1610 $D=19
M1 VSS A1 7 VSS nmos L=1.4e-07 W=7.7e-07 $X=1225 $Y=1610 $D=19
M2 Y A1 8 VSS nmos L=1.4e-07 W=7.7e-07 $X=2345 $Y=1610 $D=19
M3 8 A0 Y VSS nmos L=1.4e-07 W=7.7e-07 $X=2905 $Y=1610 $D=19
M4 VSS 6 8 VSS nmos L=1.4e-07 W=7.7e-07 $X=3465 $Y=1610 $D=19
M5 6 A0 VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=1175 $Y=4585 $D=25
M6 VDD A1 6 VDD pmos L=1.4e-07 W=1.19e-06 $X=1735 $Y=4585 $D=25
M7 9 A0 VDD VDD pmos L=1.4e-07 W=2.24e-06 $X=2365 $Y=4620 $D=25
M8 Y A1 9 VDD pmos L=1.4e-07 W=2.24e-06 $X=2855 $Y=4585 $D=25
M9 VDD 6 Y VDD pmos L=1.4e-07 W=1.19e-06 $X=3450 $Y=4620 $D=25
.ENDS
***************************************
.SUBCKT mux21 VSS VDD Y S0 A1 A0
** N=12 EP=6 IP=0 FDC=12
* PORT VSS VSS 2205 350 metal1
* PORT VDD VDD 2205 8050 metal1
* PORT Y Y 3830 3675 metal1
* PORT S0 S0 815 4935 metal1
* PORT A1 A1 1830 4305 metal1
* PORT A0 A0 2460 3675 metal1
M0 VSS S0 7 VSS nmos L=1.4e-07 W=3.5e-07 $X=850 $Y=1610 $D=19
M1 8 S0 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=1445 $Y=1190 $D=19
M2 9 A1 8 VSS nmos L=1.4e-07 W=7.7e-07 $X=1865 $Y=1190 $D=19
M3 10 A0 9 VSS nmos L=1.4e-07 W=7.7e-07 $X=2425 $Y=1190 $D=19
M4 VSS 7 10 VSS nmos L=1.4e-07 W=7.7e-07 $X=2845 $Y=1190 $D=19
M5 Y 9 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=3405 $Y=1190 $D=19
M6 VDD S0 7 VDD pmos L=1.4e-07 W=7.7e-07 $X=850 $Y=5670 $D=25
M7 11 S0 VDD VDD pmos L=1.4e-07 W=1.54e-06 $X=1445 $Y=5670 $D=25
M8 9 A0 11 VDD pmos L=1.4e-07 W=1.54e-06 $X=1865 $Y=5670 $D=25
M9 12 A1 9 VDD pmos L=1.4e-07 W=1.54e-06 $X=2425 $Y=5670 $D=25
M10 VDD 7 12 VDD pmos L=1.4e-07 W=1.54e-06 $X=2845 $Y=5670 $D=25
M11 Y 9 VDD VDD pmos L=1.4e-07 W=1.54e-06 $X=3405 $Y=5670 $D=25
.ENDS
***************************************
.SUBCKT miniALU4 Cout VSS VDD Output[3] Input1[2] Input2[2] Input1[3] Input1[1] Control[1] Output[1] Input2[1] Input2[3] Output[2] Control[0] Input1[0] Input2[0] Output[0]
** N=62 EP=17 IP=197 FDC=294
* PORT Cout Cout 29770 56035 metal2
* PORT VSS VSS -13980 22710 metal1
* PORT VDD VDD 66875 22710 metal1
* PORT Output[3] Output[3] -13980 37310 metal1
* PORT Input1[2] Input1[2] -13980 25150 metal1
* PORT Input2[2] Input2[2] -13980 20270 metal1
* PORT Input1[3] Input1[3] 16190 56035 metal2
* PORT Input1[1] Input1[1] 825 -10615 metal2
* PORT Control[1] Control[1] 46745 56035 metal2
* PORT Output[1] Output[1] 5445 -10615 metal2
* PORT Input2[1] Input2[1] 14825 -10615 metal2
* PORT Input2[3] Input2[3] 12655 56035 metal2
* PORT Output[2] Output[2] 28405 -10615 metal2
* PORT Control[0] Control[0] 32290 56035 metal2
* PORT Input1[0] Input1[0] 66875 20270 metal1
* PORT Input2[0] Input2[0] 66875 7060 metal1
* PORT Output[0] Output[0] 66875 37310 metal1
M0 VSS 4 Cout VSS nmos L=1.4e-07 W=3.5e-07 $X=30260 $Y=35245 $D=19
M1 3 49 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=30855 $Y=34825 $D=19
M2 4 Control[1] 3 VSS nmos L=1.4e-07 W=7.7e-07 $X=31275 $Y=34825 $D=19
M3 5 Control[0] 4 VSS nmos L=1.4e-07 W=7.7e-07 $X=31835 $Y=34825 $D=19
M4 VSS 52 5 VSS nmos L=1.4e-07 W=7.7e-07 $X=32255 $Y=34825 $D=19
M5 6 Input1[0] VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=32500 $Y=4995 $D=19
M6 8 53 6 VSS nmos L=1.4e-07 W=7.7e-07 $X=32920 $Y=4995 $D=19
M7 9 Control[0] 8 VSS nmos L=1.4e-07 W=1.19e-06 $X=33515 $Y=4575 $D=19
M8 10 Control[1] 9 VSS nmos L=1.4e-07 W=1.19e-06 $X=33935 $Y=4575 $D=19
M9 VSS 54 10 VSS nmos L=1.4e-07 W=1.19e-06 $X=34355 $Y=4575 $D=19
M10 11 12 VSS VSS nmos L=1.4e-07 W=3.5e-07 $X=39115 $Y=34825 $D=19
M11 VSS Control[1] 11 VSS nmos L=1.4e-07 W=3.5e-07 $X=39675 $Y=34825 $D=19
M12 12 Control[0] VSS VSS nmos L=1.4e-07 W=3.5e-07 $X=40235 $Y=34825 $D=19
M13 VDD 4 Cout VDD pmos L=1.4e-07 W=7.7e-07 $X=30120 $Y=39655 $D=25
M14 13 Control[0] VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=30715 $Y=39655 $D=25
M15 4 49 13 VDD pmos L=1.4e-07 W=1.19e-06 $X=31275 $Y=39655 $D=25
M16 13 Control[1] 4 VDD pmos L=1.4e-07 W=1.19e-06 $X=31835 $Y=39655 $D=25
M17 8 Input1[0] 14 VDD pmos L=1.4e-07 W=1.19e-06 $X=32115 $Y=9405 $D=25
M18 VDD 52 13 VDD pmos L=1.4e-07 W=1.19e-06 $X=32395 $Y=39655 $D=25
M19 14 53 8 VDD pmos L=1.4e-07 W=1.19e-06 $X=32675 $Y=9405 $D=25
M20 VDD Control[0] 14 VDD pmos L=1.4e-07 W=1.19e-06 $X=33235 $Y=9405 $D=25
M21 14 Control[1] VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=33795 $Y=9405 $D=25
M22 VDD 54 14 VDD pmos L=1.4e-07 W=1.19e-06 $X=34355 $Y=9405 $D=25
M23 15 12 11 VDD pmos L=1.4e-07 W=1.19e-06 $X=39220 $Y=39655 $D=25
M24 VDD Control[1] 15 VDD pmos L=1.4e-07 W=1.19e-06 $X=39640 $Y=39655 $D=25
M25 12 Control[0] VDD VDD pmos L=1.4e-07 W=7.7e-07 $X=40235 $Y=39655 $D=25
X26 VSS VDD 22 Input1[1] inv01 $T=20 3385 0 0 $X=20 $Y=3385
X27 VSS VDD 23 Input1[3] inv01 $T=20 18510 0 0 $X=20 $Y=18510
X28 VSS VDD Output[3] 21 inv01 $T=1980 33635 1 180 $X=20 $Y=33635
X29 VSS VDD 25 Input1[2] inv01 $T=1980 18510 0 0 $X=1980 $Y=18510
X30 VSS VDD Output[1] 30 inv01 $T=6880 3385 1 180 $X=4920 $Y=3385
X31 VSS VDD Output[2] 37 inv01 $T=26970 18510 0 0 $X=26970 $Y=18510
X32 VSS VDD 53 56 inv01 $T=37260 3385 1 180 $X=35300 $Y=3385
X33 VSS VDD 58 Input1[0] inv01 $T=41180 18510 0 0 $X=41180 $Y=18510
X34 VSS VDD 24 Control[0] inv01 $T=41180 33635 0 0 $X=41180 $Y=33635
X35 VSS VDD 52 Control[1] inv01 $T=47550 33635 1 180 $X=45590 $Y=33635
X36 VSS VDD Output[0] 61 inv01 $T=50490 33635 1 180 $X=48530 $Y=33635
X37 VDD 21 VSS Input2[3] 27 11 Input1[3] Control[1] 32 aoi222 $T=10310 33635 1 180 $X=4920 $Y=33635
X38 VDD 30 VSS Input2[1] 28 11 Input1[1] Control[1] 35 aoi222 $T=6880 3385 0 0 $X=6880 $Y=3385
X39 VDD 37 VSS Input2[2] 31 11 Input1[2] Control[1] 36 aoi222 $T=6880 18510 0 0 $X=6880 $Y=18510
X40 VDD 61 VSS Input1[0] 11 60 Input2[0] Control[1] 55 aoi222 $T=46080 18510 0 0 $X=46080 $Y=18510
X41 VSS 57 VDD Control[1] Control[0] nand02 $T=41180 18510 1 180 $X=38730 $Y=18510
X42 VSS 39 VDD Control[1] 24 nand02 $T=45590 33635 1 180 $X=43140 $Y=33635
X43 VSS VDD 28 24 22 Control[1] aoi21 $T=1980 3385 0 0 $X=1980 $Y=3385
X44 VSS VDD 27 24 23 Control[1] aoi21 $T=1980 33635 0 0 $X=1980 $Y=33635
X45 VSS VDD 31 24 25 Control[1] aoi21 $T=3940 18510 0 0 $X=3940 $Y=18510
X46 VSS VDD 60 24 58 Control[1] aoi21 $T=43140 18510 0 0 $X=43140 $Y=18510
X47 VDD VSS 38 39 Input2[3] xnor2 $T=15210 33635 1 180 $X=10310 $Y=33635
X48 VDD VSS 40 39 Input2[1] xnor2 $T=12270 3385 0 0 $X=12270 $Y=3385
X49 VDD VSS 41 39 Input2[2] xnor2 $T=12270 18510 0 0 $X=12270 $Y=18510
X50 VDD VSS 42 Input1[3] 38 xnor2 $T=15210 33635 0 0 $X=15210 $Y=33635
X51 VDD VSS 43 Input1[1] 40 xnor2 $T=17170 3385 0 0 $X=17170 $Y=3385
X52 VDD VSS 44 Input1[2] 41 xnor2 $T=17170 18510 0 0 $X=17170 $Y=18510
X53 VDD VSS 32 45 42 xnor2 $T=25010 33635 1 180 $X=20110 $Y=33635
X54 VDD VSS 35 8 43 xnor2 $T=26970 3385 1 180 $X=22070 $Y=3385
X55 VDD VSS 36 46 44 xnor2 $T=28930 18510 0 0 $X=28930 $Y=18510
X56 VDD VSS 49 39 48 xnor2 $T=38240 33635 1 180 $X=33340 $Y=33635
X57 VDD VSS 55 57 54 xnor2 $T=38730 18510 1 180 $X=33830 $Y=18510
X58 VDD VSS 54 Input1[0] 56 xnor2 $T=42160 3385 1 180 $X=37260 $Y=3385
X59 VDD VSS 56 39 Input2[0] xnor2 $T=47060 3385 1 180 $X=42160 $Y=3385
X60 VSS VDD 45 44 46 41 mux21 $T=26480 18510 1 180 $X=22070 $Y=18510
X61 VSS VDD 48 42 45 38 mux21 $T=25010 33635 0 0 $X=25010 $Y=33635
X62 VSS VDD 46 43 8 40 mux21 $T=26970 3385 0 0 $X=26970 $Y=3385
.ENDS
***************************************
