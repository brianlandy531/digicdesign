* SPICE NETLIST
***************************************

.SUBCKT mimcap_g13 plus minus
.ENDS
***************************************
.SUBCKT spiral_inductor_lvs pos neg
.ENDS
***************************************
.SUBCKT inv01 VSS VDD Y A
** N=4 EP=4 IP=0 FDC=2
* PORT VSS VSS 980 350 metal1
* PORT VDD VDD 980 8050 metal1
* PORT Y Y 1435 3675 metal1
* PORT A A 805 3675 metal1
M0 Y A VSS VSS nmos L=1.4e-07 W=3.5e-07 $X=910 $Y=1820 $D=19
M1 Y A VDD VDD pmos L=1.4e-07 W=7.7e-07 $X=910 $Y=5600 $D=25
.ENDS
***************************************
.SUBCKT xnor2 VDD VSS Y A0 A1
** N=9 EP=5 IP=0 FDC=10
* PORT VDD VDD 2450 8050 metal1
* PORT VSS VSS 2450 350 metal1
* PORT Y Y 3955 3675 metal1
* PORT A0 A0 980 3675 metal1
* PORT A1 A1 2555 3675 metal1
M0 7 A0 6 VSS nmos L=1.4e-07 W=7.7e-07 $X=805 $Y=1610 $D=19
M1 VSS A1 7 VSS nmos L=1.4e-07 W=7.7e-07 $X=1225 $Y=1610 $D=19
M2 Y A1 8 VSS nmos L=1.4e-07 W=7.7e-07 $X=2345 $Y=1610 $D=19
M3 8 A0 Y VSS nmos L=1.4e-07 W=7.7e-07 $X=2905 $Y=1610 $D=19
M4 VSS 6 8 VSS nmos L=1.4e-07 W=7.7e-07 $X=3465 $Y=1610 $D=19
M5 6 A0 VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=1175 $Y=4585 $D=25
M6 VDD A1 6 VDD pmos L=1.4e-07 W=1.19e-06 $X=1735 $Y=4585 $D=25
M7 9 A0 VDD VDD pmos L=1.4e-07 W=2.24e-06 $X=2365 $Y=4620 $D=25
M8 Y A1 9 VDD pmos L=1.4e-07 W=2.24e-06 $X=2855 $Y=4585 $D=25
M9 VDD 6 Y VDD pmos L=1.4e-07 W=1.19e-06 $X=3450 $Y=4620 $D=25
.ENDS
***************************************
.SUBCKT oai222 VDD Y VSS A0 A1 B1 B0 C0 C1
** N=14 EP=9 IP=0 FDC=12
* PORT VDD VDD 2695 8050 metal1
* PORT Y Y 1855 3675 metal1
* PORT VSS VSS 2695 350 metal1
* PORT A0 A0 595 3675 metal1
* PORT A1 A1 1225 3675 metal1
* PORT B1 B1 2485 3675 metal1
* PORT B0 B0 3115 3675 metal1
* PORT C0 C0 3745 3675 metal1
* PORT C1 C1 4375 3675 metal1
M0 Y A0 10 VSS nmos L=1.4e-07 W=1.19e-06 $X=805 $Y=1610 $D=19
M1 10 A1 Y VSS nmos L=1.4e-07 W=1.19e-06 $X=1365 $Y=1610 $D=19
M2 10 B1 11 VSS nmos L=1.4e-07 W=1.19e-06 $X=2485 $Y=1610 $D=19
M3 11 B0 10 VSS nmos L=1.4e-07 W=1.19e-06 $X=3045 $Y=1610 $D=19
M4 VSS C0 11 VSS nmos L=1.4e-07 W=1.19e-06 $X=3605 $Y=1610 $D=19
M5 11 C1 VSS VSS nmos L=1.4e-07 W=1.19e-06 $X=4165 $Y=1610 $D=19
M6 12 A0 VDD VDD pmos L=1.4e-07 W=2.52e-06 $X=1365 $Y=4690 $D=25
M7 Y A1 12 VDD pmos L=1.4e-07 W=2.52e-06 $X=1785 $Y=4690 $D=25
M8 13 B1 Y VDD pmos L=1.4e-07 W=2.52e-06 $X=2345 $Y=4690 $D=25
M9 VDD B0 13 VDD pmos L=1.4e-07 W=2.52e-06 $X=2765 $Y=4690 $D=25
M10 14 C0 VDD VDD pmos L=1.4e-07 W=2.52e-06 $X=3325 $Y=4690 $D=25
M11 Y C1 14 VDD pmos L=1.4e-07 W=2.52e-06 $X=3745 $Y=4690 $D=25
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=13 FDC=14
X0 2 3 4 1 inv01 $T=7350 0 1 180 $X=5390 $Y=0
X1 3 6 2 5 7 8 9 10 11 oai222 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT aoi21 VSS VDD Y A1 A0 B0
** N=8 EP=6 IP=0 FDC=6
* PORT VSS VSS 1470 350 metal1
* PORT VDD VDD 1470 8050 metal1
* PORT Y Y 2485 3675 metal1
* PORT A1 A1 560 3675 metal1
* PORT A0 A0 1190 3045 metal1
* PORT B0 B0 1855 4305 metal1
M0 7 A1 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=805 $Y=1170 $D=19
M1 Y A0 7 VSS nmos L=1.4e-07 W=7.7e-07 $X=1225 $Y=1170 $D=19
M2 VSS B0 Y VSS nmos L=1.4e-07 W=3.5e-07 $X=1820 $Y=1590 $D=19
M3 VDD A1 8 VDD pmos L=1.4e-07 W=1.19e-06 $X=805 $Y=6020 $D=25
M4 8 A0 VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=1365 $Y=6020 $D=25
M5 Y B0 8 VDD pmos L=1.4e-07 W=1.19e-06 $X=1925 $Y=6020 $D=25
.ENDS
***************************************
.SUBCKT xor2 VSS VDD Y A1 A0
** N=10 EP=5 IP=0 FDC=12
* PORT VSS VSS 2450 350 metal1
* PORT VDD VDD 2450 8050 metal1
* PORT Y Y 4445 3150 metal1
* PORT A1 A1 2555 3150 metal1
* PORT A0 A0 840 3150 metal1
M0 7 A0 6 VSS nmos L=1.4e-07 W=7.7e-07 $X=805 $Y=1330 $D=19
M1 VSS A1 7 VSS nmos L=1.4e-07 W=7.7e-07 $X=1225 $Y=1330 $D=19
M2 8 6 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=1785 $Y=1330 $D=19
M3 9 A1 8 VSS nmos L=1.4e-07 W=7.7e-07 $X=2345 $Y=1330 $D=19
M4 8 A0 9 VSS nmos L=1.4e-07 W=7.7e-07 $X=2905 $Y=1330 $D=19
M5 Y 9 VSS VSS nmos L=1.4e-07 W=3.5e-07 $X=4025 $Y=1330 $D=19
M6 6 A0 VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=875 $Y=5880 $D=25
M7 VDD A1 6 VDD pmos L=1.4e-07 W=1.19e-06 $X=1435 $Y=5880 $D=25
M8 9 6 VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=1995 $Y=5880 $D=25
M9 10 A1 9 VDD pmos L=1.4e-07 W=2.24e-06 $X=2590 $Y=4830 $D=25
M10 VDD A0 10 VDD pmos L=1.4e-07 W=2.24e-06 $X=3010 $Y=4830 $D=25
M11 Y 9 VDD VDD pmos L=1.4e-07 W=7.7e-07 $X=3605 $Y=4830 $D=25
.ENDS
***************************************
.SUBCKT mux21 VSS VDD Y S0 A1 A0
** N=12 EP=6 IP=0 FDC=12
* PORT VSS VSS 2205 350 metal1
* PORT VDD VDD 2205 8050 metal1
* PORT Y Y 3830 3675 metal1
* PORT S0 S0 815 4935 metal1
* PORT A1 A1 1830 4305 metal1
* PORT A0 A0 2460 3675 metal1
M0 VSS S0 7 VSS nmos L=1.4e-07 W=3.5e-07 $X=850 $Y=1610 $D=19
M1 8 S0 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=1445 $Y=1190 $D=19
M2 9 A1 8 VSS nmos L=1.4e-07 W=7.7e-07 $X=1865 $Y=1190 $D=19
M3 10 A0 9 VSS nmos L=1.4e-07 W=7.7e-07 $X=2425 $Y=1190 $D=19
M4 VSS 7 10 VSS nmos L=1.4e-07 W=7.7e-07 $X=2845 $Y=1190 $D=19
M5 Y 9 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=3405 $Y=1190 $D=19
M6 VDD S0 7 VDD pmos L=1.4e-07 W=7.7e-07 $X=850 $Y=5670 $D=25
M7 11 S0 VDD VDD pmos L=1.4e-07 W=1.54e-06 $X=1445 $Y=5670 $D=25
M8 9 A0 11 VDD pmos L=1.4e-07 W=1.54e-06 $X=1865 $Y=5670 $D=25
M9 12 A1 9 VDD pmos L=1.4e-07 W=1.54e-06 $X=2425 $Y=5670 $D=25
M10 VDD 7 12 VDD pmos L=1.4e-07 W=1.54e-06 $X=2845 $Y=5670 $D=25
M11 Y 9 VDD VDD pmos L=1.4e-07 W=1.54e-06 $X=3405 $Y=5670 $D=25
.ENDS
***************************************
.SUBCKT inv02 VSS VDD Y A
** N=4 EP=4 IP=0 FDC=2
* PORT VSS VSS 980 350 metal1
* PORT VDD VDD 980 8050 metal1
* PORT Y Y 1330 3675 metal1
* PORT A A 700 3675 metal1
M0 Y A VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=805 $Y=1750 $D=19
M1 Y A VDD VDD pmos L=1.4e-07 W=1.54e-06 $X=805 $Y=4970 $D=25
.ENDS
***************************************
.SUBCKT nand02 VSS Y VDD A1 A0
** N=6 EP=5 IP=0 FDC=4
* PORT VSS VSS 1225 350 metal1
* PORT Y Y 1925 3675 metal1
* PORT VDD VDD 1225 8050 metal1
* PORT A1 A1 665 3675 metal1
* PORT A0 A0 1295 4305 metal1
M0 6 A1 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=875 $Y=1190 $D=19
M1 Y A0 6 VSS nmos L=1.4e-07 W=7.7e-07 $X=1295 $Y=1190 $D=19
M2 Y A1 VDD VDD pmos L=1.4e-07 W=1.05e-06 $X=875 $Y=6160 $D=25
M3 VDD A0 Y VDD pmos L=1.4e-07 W=1.05e-06 $X=1435 $Y=6160 $D=25
.ENDS
***************************************
.SUBCKT buf02 VSS VDD Y A
** N=5 EP=4 IP=0 FDC=4
* PORT VSS VSS 1225 350 metal1
* PORT VDD VDD 1225 8050 metal1
* PORT Y Y 1875 3675 metal1
* PORT A A 720 3675 metal1
M0 VSS A 5 VSS nmos L=1.4e-07 W=3.5e-07 $X=860 $Y=1610 $D=19
M1 Y 5 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=1455 $Y=1190 $D=19
M2 VDD A 5 VDD pmos L=1.4e-07 W=7.7e-07 $X=860 $Y=5670 $D=25
M3 Y 5 VDD VDD pmos L=1.4e-07 W=1.54e-06 $X=1455 $Y=5670 $D=25
.ENDS
***************************************
.SUBCKT miniALU16 VSS VDD Cout Input2[7] Input2[8] Input1[2] Output[2] Output[8] Input2[2] Input1[1] Input1[13] Input1[8] Input1[7] Input2[13] Output[7] Output[1] Input2[10] Output[13] Input2[1] Input1[10]
+ Output[10] Input1[9] Input2[4] Output[9] Input2[9] Input2[3] Input1[3] Input1[12] Output[3] Input1[4] Input2[12] Control[0] Output[4] Input1[11] Control[1] Input2[0] Output[12] Input2[5] Output[0] Input1[0]
+ Input1[15] Input1[6] Input2[11] Input2[6] Input1[14] Output[15] Input1[5] Input2[14] Output[14] Output[5] Output[6] Input2[15] Output[11]
** N=191 EP=53 IP=729 FDC=1116
* PORT VSS VSS -27980 45400 metal1
* PORT VDD VDD 121940 45400 metal1
* PORT Cout Cout 60430 -24615 metal2
* PORT Input2[7] Input2[7] -27980 37310 metal1
* PORT Input2[8] Input2[8] -27980 56775 metal1
* PORT Input1[2] Input1[2] -27980 69460 metal1
* PORT Output[2] Output[2] -27980 67020 metal1
* PORT Output[8] Output[8] -27980 51895 metal1
* PORT Input2[2] Input2[2] -27980 54335 metal1
* PORT Input1[1] Input1[1] -27980 82055 metal1
* PORT Input1[13] Input1[13] -27980 21555 metal1
* PORT Input1[8] Input1[8] -27980 39750 metal1
* PORT Input1[7] Input1[7] -27980 6430 metal1
* PORT Input2[13] Input2[13] 16165 -24615 metal2
* PORT Output[7] Output[7] 10765 -24615 metal2
* PORT Output[1] Output[1] 6425 115410 metal2
* PORT Input2[10] Input2[10] 38625 -24615 metal2
* PORT Output[13] Output[13] 18605 -24615 metal2
* PORT Input2[1] Input2[1] 14615 115410 metal2
* PORT Input1[10] Input1[10] 26270 -24615 metal2
* PORT Output[10] Output[10] 23015 -24615 metal2
* PORT Input1[9] Input1[9] 37960 115410 metal2
* PORT Input2[4] Input2[4] 31765 -24615 metal2
* PORT Output[9] Output[9] 41215 115410 metal2
* PORT Input2[9] Input2[9] 34215 115410 metal2
* PORT Input2[3] Input2[3] 44750 -24615 metal2
* PORT Input1[3] Input1[3] 44820 115410 metal2
* PORT Input1[12] Input1[12] 84300 115410 metal2
* PORT Output[3] Output[3] 48075 115410 metal2
* PORT Input1[4] Input1[4] 55075 -24615 metal2
* PORT Input2[12] Input2[12] 80975 115410 metal2
* PORT Control[0] Control[0] 35615 -24615 metal2
* PORT Output[4] Output[4] 50035 -24615 metal2
* PORT Input1[11] Input1[11] 121940 54875 metal1
* PORT Control[1] Control[1] 57210 115410 metal2
* PORT Input2[0] Input2[0] 51575 115410 metal2
* PORT Output[12] Output[12] 74955 115410 metal2
* PORT Input2[5] Input2[5] 63335 -24615 metal2
* PORT Output[0] Output[0] 62705 115410 metal2
* PORT Input1[0] Input1[0] 65365 115410 metal2
* PORT Input1[15] Input1[15] 121940 65120 metal1
* PORT Input1[6] Input1[6] 121940 28965 metal1
* PORT Input2[11] Input2[11] 121940 52435 metal1
* PORT Input2[6] Input2[6] 121940 24085 metal1
* PORT Input1[14] Input1[14] 121940 41650 metal1
* PORT Output[15] Output[15] 69635 115410 metal2
* PORT Input1[5] Input1[5] 121940 6430 metal1
* PORT Input2[14] Input2[14] 121940 26525 metal1
* PORT Output[14] Output[14] 121940 36770 metal1
* PORT Output[5] Output[5] 86295 -24615 metal2
* PORT Output[6] Output[6] 121940 21645 metal1
* PORT Input2[15] Input2[15] 121940 67560 metal1
* PORT Output[11] Output[11] 121940 39210 metal1
M0 VSS Control[0] 1 VSS nmos L=1.4e-07 W=3.5e-07 $X=56685 $Y=65075 $D=19
M1 4 Control[1] VSS VSS nmos L=1.4e-07 W=3.5e-07 $X=57245 $Y=19700 $D=19
M2 5 Control[1] VSS VSS nmos L=1.4e-07 W=3.5e-07 $X=57245 $Y=65075 $D=19
M3 VSS Control[0] 4 VSS nmos L=1.4e-07 W=3.5e-07 $X=57805 $Y=19700 $D=19
M4 VSS 1 5 VSS nmos L=1.4e-07 W=3.5e-07 $X=57805 $Y=65075 $D=19
M5 6 45 VSS VSS nmos L=1.4e-07 W=7.7e-07 $X=59275 $Y=34825 $D=19
M6 7 Control[0] 6 VSS nmos L=1.4e-07 W=7.7e-07 $X=59695 $Y=34825 $D=19
M7 8 Control[1] 7 VSS nmos L=1.4e-07 W=7.7e-07 $X=60255 $Y=34825 $D=19
M8 VSS 138 8 VSS nmos L=1.4e-07 W=7.7e-07 $X=60675 $Y=34825 $D=19
M9 Cout 7 VSS VSS nmos L=1.4e-07 W=3.5e-07 $X=61270 $Y=35245 $D=19
M10 10 137 VSS VSS nmos L=1.4e-07 W=1.19e-06 $X=63545 $Y=49950 $D=19
M11 11 Control[1] 10 VSS nmos L=1.4e-07 W=1.19e-06 $X=63965 $Y=49950 $D=19
M12 12 Control[0] 11 VSS nmos L=1.4e-07 W=1.19e-06 $X=64385 $Y=49950 $D=19
M13 13 149 12 VSS nmos L=1.4e-07 W=7.7e-07 $X=64980 $Y=50370 $D=19
M14 VSS Input1[0] 13 VSS nmos L=1.4e-07 W=7.7e-07 $X=65400 $Y=50370 $D=19
M15 VDD Control[0] 1 VDD pmos L=1.4e-07 W=7.7e-07 $X=56685 $Y=69905 $D=25
M16 14 Control[1] 4 VDD pmos L=1.4e-07 W=1.19e-06 $X=57245 $Y=24530 $D=25
M17 15 Control[1] VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=57280 $Y=69905 $D=25
M18 VDD Control[0] 14 VDD pmos L=1.4e-07 W=1.19e-06 $X=57665 $Y=24530 $D=25
M19 5 1 15 VDD pmos L=1.4e-07 W=1.19e-06 $X=57700 $Y=69905 $D=25
M20 16 45 VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=59135 $Y=39655 $D=25
M21 7 Control[1] 16 VDD pmos L=1.4e-07 W=1.19e-06 $X=59695 $Y=39655 $D=25
M22 16 138 7 VDD pmos L=1.4e-07 W=1.19e-06 $X=60255 $Y=39655 $D=25
M23 VDD Control[0] 16 VDD pmos L=1.4e-07 W=1.19e-06 $X=60815 $Y=39655 $D=25
M24 Cout 7 VDD VDD pmos L=1.4e-07 W=7.7e-07 $X=61410 $Y=39655 $D=25
M25 17 137 VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=63545 $Y=54780 $D=25
M26 VDD Control[1] 17 VDD pmos L=1.4e-07 W=1.19e-06 $X=64105 $Y=54780 $D=25
M27 17 Control[0] VDD VDD pmos L=1.4e-07 W=1.19e-06 $X=64665 $Y=54780 $D=25
M28 12 149 17 VDD pmos L=1.4e-07 W=1.19e-06 $X=65225 $Y=54780 $D=25
M29 17 Input1[0] 12 VDD pmos L=1.4e-07 W=1.19e-06 $X=65785 $Y=54780 $D=25
X30 VSS VDD 29 Input2[8] inv01 $T=20 48760 0 0 $X=20 $Y=48760
X31 VSS VDD 30 Input2[2] inv01 $T=20 79010 0 0 $X=20 $Y=79010
X32 VSS VDD 35 Input1[8] inv01 $T=1980 48760 0 0 $X=1980 $Y=48760
X33 VSS VDD 36 Input1[2] inv01 $T=1980 79010 0 0 $X=1980 $Y=79010
X34 VSS VDD 41 Input2[7] inv01 $T=4920 18510 0 0 $X=4920 $Y=18510
X35 VSS VDD 56 Input2[13] inv01 $T=11780 18510 0 0 $X=11780 $Y=18510
X36 VSS VDD 59 Input1[13] inv01 $T=12270 33635 0 0 $X=12270 $Y=33635
X37 VSS VDD 73 Input2[10] inv01 $T=20110 3385 0 0 $X=20110 $Y=3385
X38 VSS VDD 68 Input1[1] inv01 $T=24520 79010 1 180 $X=22560 $Y=79010
X39 VSS VDD 88 Input1[9] inv01 $T=27460 79010 0 0 $X=27460 $Y=79010
X40 VSS VDD 104 Input2[4] inv01 $T=37260 3385 0 0 $X=37260 $Y=3385
X41 VSS VDD 114 Input2[3] inv01 $T=45100 18510 0 0 $X=45100 $Y=18510
X42 VSS VDD 125 Control[0] inv01 $T=49510 18510 0 0 $X=49510 $Y=18510
X43 VSS VDD 45 Control[1] inv01 $T=53430 79010 1 180 $X=51470 $Y=79010
X44 VSS VDD 69 Control[1] inv01 $T=51960 63885 0 0 $X=51960 $Y=63885
X45 VSS VDD 133 Input2[0] inv01 $T=53920 63885 0 0 $X=53920 $Y=63885
X46 VSS VDD 135 Input2[12] inv01 $T=65680 79010 1 180 $X=63720 $Y=79010
X47 VSS VDD 49 154 inv01 $T=67640 79010 1 180 $X=65680 $Y=79010
X48 VSS VDD 149 131 inv01 $T=68620 48760 1 180 $X=66660 $Y=48760
X49 VSS VDD 155 154 inv01 $T=67640 79010 0 0 $X=67640 $Y=79010
X50 VSS VDD 163 Input1[15] inv01 $T=72540 79010 0 0 $X=72540 $Y=79010
X51 VSS VDD 176 Input2[5] inv01 $T=78910 3385 0 0 $X=78910 $Y=3385
X52 VSS VDD 166 Input2[15] inv01 $T=86750 79010 1 180 $X=84790 $Y=79010
X53 VSS VDD 179 Input2[14] inv01 $T=89690 33635 1 180 $X=87730 $Y=33635
X54 VSS VDD 184 Input1[6] inv01 $T=90670 18510 1 180 $X=88710 $Y=18510
X55 VSS VDD 190 Input1[11] inv01 $T=93120 48760 1 180 $X=91160 $Y=48760
X56 VDD VSS 33 Input1[7] 31 xnor2 $T=20 3385 0 0 $X=20 $Y=3385
X57 VDD VSS 31 28 Input2[7] xnor2 $T=20 18510 0 0 $X=20 $Y=18510
X58 VDD VSS 40 28 Input2[8] xnor2 $T=20 33635 0 0 $X=20 $Y=33635
X59 VDD VSS 34 Input1[2] 32 xnor2 $T=20 63885 0 0 $X=20 $Y=63885
X60 VDD VSS 53 28 Input2[13] xnor2 $T=6880 18510 0 0 $X=6880 $Y=18510
X61 VDD VSS 63 Input1[8] 40 xnor2 $T=12270 48760 0 0 $X=12270 $Y=48760
X62 VDD VSS 64 28 Input2[10] xnor2 $T=13740 18510 0 0 $X=13740 $Y=18510
X63 VDD VSS 32 70 Input2[2] xnor2 $T=19130 63885 1 180 $X=14230 $Y=63885
X64 VDD VSS 71 Input1[10] 64 xnor2 $T=23540 18510 1 180 $X=18640 $Y=18510
X65 VDD VSS 76 70 Input2[1] xnor2 $T=19130 63885 0 0 $X=19130 $Y=63885
X66 VDD VSS 78 Input1[13] 53 xnor2 $T=19620 33635 0 0 $X=19620 $Y=33635
X67 VDD VSS 86 Input1[1] 76 xnor2 $T=24030 63885 0 0 $X=24030 $Y=63885
X68 VDD VSS 102 70 Input2[4] xnor2 $T=32360 3385 0 0 $X=32360 $Y=3385
X69 VDD VSS 99 70 Input2[3] xnor2 $T=32850 18510 0 0 $X=32850 $Y=18510
X70 VDD VSS 87 Input1[9] 98 xnor2 $T=35790 48760 0 0 $X=35790 $Y=48760
X71 VDD VSS 92 Input1[3] 99 xnor2 $T=43140 33635 1 180 $X=38240 $Y=33635
X72 VDD VSS 98 28 Input2[9] xnor2 $T=45590 48760 1 180 $X=40690 $Y=48760
X73 VDD VSS 103 Input1[12] 108 xnor2 $T=46570 79010 1 180 $X=41670 $Y=79010
X74 VDD VSS 109 Input1[4] 102 xnor2 $T=48530 3385 1 180 $X=43630 $Y=3385
X75 VDD VSS 108 28 Input2[12] xnor2 $T=46570 79010 0 0 $X=46570 $Y=79010
X76 VDD VSS 112 Input1[11] 113 xnor2 $T=51960 63885 1 180 $X=47060 $Y=63885
X77 VDD VSS 131 70 Input2[0] xnor2 $T=50490 48760 0 0 $X=50490 $Y=48760
X78 VDD VSS 146 70 Input2[5] xnor2 $T=59800 3385 0 0 $X=59800 $Y=3385
X79 VDD VSS 138 28 148 xnor2 $T=67640 33635 1 180 $X=62740 $Y=33635
X80 VDD VSS 142 Input1[6] 144 xnor2 $T=73520 18510 1 180 $X=68620 $Y=18510
X81 VDD VSS 137 Input1[0] 131 xnor2 $T=68620 48760 0 0 $X=68620 $Y=48760
X82 VDD VSS 156 Input1[14] 162 xnor2 $T=77440 33635 1 180 $X=72540 $Y=33635
X83 VDD VSS 113 28 Input2[11] xnor2 $T=77930 63885 1 180 $X=73030 $Y=63885
X84 VDD VSS 144 28 Input2[6] xnor2 $T=73520 18510 0 0 $X=73520 $Y=18510
X85 VDD VSS 153 Input1[5] 146 xnor2 $T=78910 3385 1 180 $X=74010 $Y=3385
X86 VDD VSS 162 28 Input2[14] xnor2 $T=77930 48760 0 0 $X=77930 $Y=48760
X87 VDD VSS 173 28 Input2[15] xnor2 $T=85280 63885 0 0 $X=85280 $Y=63885
X88 VDD VSS 177 Input1[15] 173 xnor2 $T=91650 79010 1 180 $X=86750 $Y=79010
X89 VDD Output[8] VSS 45 44 42 29 35 37 oai222 $T=9330 48760 1 180 $X=3940 $Y=48760
X90 VDD Output[2] VSS 45 38 43 30 36 37 oai222 $T=9330 79010 1 180 $X=3940 $Y=79010
X91 VDD Output[13] VSS 69 66 54 56 59 37 oai222 $T=19620 33635 1 180 $X=14230 $Y=33635
X92 VDD Output[15] VSS 69 171 159 166 163 154 oai222 $T=79890 79010 1 180 $X=74500 $Y=79010
X93 Input1[7] VSS VDD 55 45 Output[7] 51 52 41 55 37 ICV_1 $T=9820 3385 0 0 $X=9820 $Y=3385
X94 Input2[1] VSS VDD 65 45 Output[1] 61 58 65 68 37 ICV_1 $T=15210 79010 0 0 $X=15210 $Y=79010
X95 Input1[10] VSS VDD 80 45 Output[10] 77 79 73 80 37 ICV_1 $T=22070 3385 0 0 $X=22070 $Y=3385
X96 Input2[9] VSS VDD 90 45 Output[9] 89 83 90 88 37 ICV_1 $T=29420 79010 0 0 $X=29420 $Y=79010
X97 Input1[3] VSS VDD 126 45 Output[3] 115 122 114 126 37 ICV_1 $T=48040 33635 0 0 $X=48040 $Y=33635
X98 Input1[4] VSS VDD 129 45 Output[4] 110 127 104 129 37 ICV_1 $T=49510 3385 0 0 $X=49510 $Y=3385
X99 Input1[12] VSS VDD 136 69 Output[12] 106 132 135 136 37 ICV_1 $T=56370 79010 0 0 $X=56370 $Y=79010
X100 Input1[0] VSS VDD 147 45 Output[0] 141 37 147 133 151 ICV_1 $T=60780 63885 0 0 $X=60780 $Y=63885
X101 Input1[14] VSS VDD 180 69 Output[14] 158 172 179 180 37 ICV_1 $T=80380 33635 0 0 $X=80380 $Y=33635
X102 Input2[6] VSS VDD 181 45 Output[6] 152 175 181 184 37 ICV_1 $T=81360 18510 0 0 $X=81360 $Y=18510
X103 Input1[5] VSS VDD 189 45 Output[5] 161 178 176 189 37 ICV_1 $T=83810 3385 0 0 $X=83810 $Y=3385
X104 Input2[11] VSS VDD 188 69 Output[11] 120 185 188 190 37 ICV_1 $T=83810 48760 0 0 $X=83810 $Y=48760
X105 VSS VDD 54 4 Input1[13] 49 aoi21 $T=12270 33635 1 180 $X=9330 $Y=33635
X106 VSS VDD 42 4 Input1[8] 49 aoi21 $T=12270 48760 1 180 $X=9330 $Y=48760
X107 VSS VDD 43 4 Input1[2] 49 aoi21 $T=12270 79010 1 180 $X=9330 $Y=79010
X108 VSS VDD 58 4 Input1[1] 49 aoi21 $T=12270 79010 0 0 $X=12270 $Y=79010
X109 VSS VDD 52 4 Input1[7] 49 aoi21 $T=20110 3385 1 180 $X=17170 $Y=3385
X110 VSS VDD 83 4 Input1[9] 49 aoi21 $T=24520 79010 0 0 $X=24520 $Y=79010
X111 VSS VDD 79 4 Input1[10] 49 aoi21 $T=32360 3385 1 180 $X=29420 $Y=3385
X112 VSS VDD 132 4 Input1[12] 49 aoi21 $T=53430 79010 0 0 $X=53430 $Y=79010
X113 VSS VDD 122 4 Input1[3] 49 aoi21 $T=58330 33635 1 180 $X=55390 $Y=33635
X114 VSS VDD 127 4 Input1[4] 49 aoi21 $T=56860 3385 0 0 $X=56860 $Y=3385
X115 VSS VDD 151 4 Input1[0] 49 aoi21 $T=71070 63885 1 180 $X=68130 $Y=63885
X116 VSS VDD 159 4 Input1[15] 155 aoi21 $T=69600 79010 0 0 $X=69600 $Y=79010
X117 VSS VDD 172 4 Input1[14] 49 aoi21 $T=77440 33635 0 0 $X=77440 $Y=33635
X118 VSS VDD 175 4 Input1[6] 49 aoi21 $T=78420 18510 0 0 $X=78420 $Y=18510
X119 VSS VDD 178 4 Input1[5] 49 aoi21 $T=80870 3385 0 0 $X=80870 $Y=3385
X120 VSS VDD 185 4 Input1[11] 49 aoi21 $T=82340 63885 0 0 $X=82340 $Y=63885
X121 VSS VDD 51 33 39 xor2 $T=4920 3385 0 0 $X=4920 $Y=3385
X122 VSS VDD 38 34 46 xor2 $T=9820 63885 1 180 $X=4920 $Y=63885
X123 VSS VDD 44 63 47 xor2 $T=22070 48760 1 180 $X=17170 $Y=48760
X124 VSS VDD 77 71 84 xor2 $T=28440 18510 1 180 $X=23540 $Y=18510
X125 VSS VDD 66 78 85 xor2 $T=29420 33635 1 180 $X=24520 $Y=33635
X126 VSS VDD 89 87 82 xor2 $T=26480 48760 0 0 $X=26480 $Y=48760
X127 VSS VDD 61 86 12 xor2 $T=38240 63885 1 180 $X=33340 $Y=63885
X128 VSS VDD 106 103 100 xor2 $T=36770 79010 0 0 $X=36770 $Y=79010
X129 VSS VDD 110 109 101 xor2 $T=40200 18510 0 0 $X=40200 $Y=18510
X130 VSS VDD 115 92 57 xor2 $T=43140 33635 0 0 $X=43140 $Y=33635
X131 VSS VDD 120 112 91 xor2 $T=45590 48760 0 0 $X=45590 $Y=48760
X132 VSS VDD 141 137 134 xor2 $T=57840 48760 0 0 $X=57840 $Y=48760
X133 VSS VDD 152 142 139 xor2 $T=63720 18510 0 0 $X=63720 $Y=18510
X134 VSS VDD 158 156 95 xor2 $T=67640 33635 0 0 $X=67640 $Y=33635
X135 VSS VDD 161 153 105 xor2 $T=69110 3385 0 0 $X=69110 $Y=3385
X136 VSS VDD 171 177 170 xor2 $T=84790 79010 1 180 $X=79890 $Y=79010
X137 VSS VDD 47 33 39 31 mux21 $T=4920 33635 0 0 $X=4920 $Y=33635
X138 VSS VDD 57 34 46 32 mux21 $T=9820 63885 0 0 $X=9820 $Y=63885
X139 VSS VDD 82 63 47 40 mux21 $T=22070 48760 0 0 $X=22070 $Y=48760
X140 VSS VDD 91 71 84 64 mux21 $T=28440 18510 0 0 $X=28440 $Y=18510
X141 VSS VDD 46 86 12 76 mux21 $T=33340 63885 1 180 $X=28930 $Y=63885
X142 VSS VDD 95 78 85 53 mux21 $T=29420 33635 0 0 $X=29420 $Y=33635
X143 VSS VDD 84 87 82 98 mux21 $T=35790 48760 1 180 $X=31380 $Y=48760
X144 VSS VDD 101 92 57 99 mux21 $T=33830 33635 0 0 $X=33830 $Y=33635
X145 VSS VDD 85 103 100 108 mux21 $T=42650 63885 1 180 $X=38240 $Y=63885
X146 VSS VDD 105 109 101 102 mux21 $T=43630 3385 1 180 $X=39220 $Y=3385
X147 VSS VDD 100 112 91 113 mux21 $T=47060 63885 1 180 $X=42650 $Y=63885
X148 VSS VDD 39 142 139 144 mux21 $T=63720 18510 1 180 $X=59310 $Y=18510
X149 VSS VDD 139 153 105 146 mux21 $T=69110 3385 1 180 $X=64700 $Y=3385
X150 VSS VDD 170 156 95 162 mux21 $T=73520 48760 0 0 $X=73520 $Y=48760
X151 VSS VDD 148 177 170 173 mux21 $T=82340 63885 1 180 $X=77930 $Y=63885
X152 VSS VDD 37 5 inv02 $T=58820 63885 0 0 $X=58820 $Y=63885
X153 VSS VDD 154 5 inv02 $T=71070 63885 0 0 $X=71070 $Y=63885
X154 VSS 117 VDD Control[1] 125 nand02 $T=53920 18510 1 180 $X=51470 $Y=18510
X155 VSS 134 VDD Control[1] Control[0] nand02 $T=57840 48760 1 180 $X=55390 $Y=48760
X156 VSS VDD 28 117 buf02 $T=49510 18510 1 180 $X=47060 $Y=18510
X157 VSS VDD 70 117 buf02 $T=56370 18510 1 180 $X=53920 $Y=18510
.ENDS
***************************************
