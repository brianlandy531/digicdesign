* Example circuit file for simulating PEX

.INCLUDE "/home/bxl1703/Pyxis_SPT_HEP/ic_projects/Pyxis_SPT/digicdesign/inv2/inv2.cal/inv2.pex.netlist"

.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_33
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_lwt
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_hwt
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_BIP
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_BIP_NPN
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo DIO
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo DIO_33
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_RES
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo MOS_CAP
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/res.spi res_t











* - Instantiate your parasitic netlist and add the load capacitor
** FORMAT : 
* XLAYOUT [all inputs as listed by the ".subckt" line in the included netlist, in the order that they appear there] [name of the subcircuit as listed in the included netlist]
XLAYOUT GROUND VOUT VIN INV2
COUT VOUT 0 120f

* - Analysis Setup - DC sweep
* FORMAT : .DC [name] [low] [high] [step]
.DC VFORCE__VIN 0 1.20 0.01

* - Analysis Setup - Trans
* FORMAT : .TRAN [start time] [end time] [time step]
.TRAN 0 20n 0.001n

* --- Forces
* FORMAT -- PULSE : [name] [port] [reference (0 means ground)] PULSE [low] [high] [delay] [fall time] [rise time] [pulse width] [period]
*
* FORMAT -- DC    : [name] [port] [reference (0 means ground)] DC [voltage]
*
VFORCE__Vin VIN 0 PULSE (0 1.2 5n 0.1n 0.1n 5n 10n)
VFORCE__Vdd VDD 0 DC 1.2
*VFORCE__VSS VSS 0 DC 0

VFORCE__GROUND GROUND 0 DC 0

* --- Waveform Outputs
.PLOT DC V(VIN)
.PLOT DC V(VOUT)
.PLOT TRAN V(VIN)
.PLOT TRAN V(VOUT)

* --- Params
.TEMP 25

