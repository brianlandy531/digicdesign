* Component: $PYXIS_SPT/digicdesign/4bitripplecarry Viewpoint: prelayout

.INCLUDE "$PYXIS_SPT/digicdesign/4bitripplecarry/prelayout/netlist.spi"
.INCLUDE "$GENERIC13/models/include_all"
.OPTION AEX
.OPTION ENGNOT
.OPTION LIMPROBE=10000.0
.OPTION NOASCII

* - Analysis Setup - DCOP
.OPTION PROBEOP2
.OP

* - Analysis Setup - Trans
.TRAN 0 1000n

* --- Forces
VFORCE__VDD VDD GROUND DC 1.08
VFORCE___ground GROUND GROUND DC 0
VFORCE__Cin0 CIN0 GROUND PATTERN 1.08 0 0 .01n .01n 20n 101 R=-1
VFORCE__B0 B0 GROUND PATTERN 1.08 0 0 .01n .01n 20n 011 R=-1
VFORCE__B1 B1 GROUND PATTERN 1.08 0 0 .01n .01n 20n 010 R=-1
VFORCE__B2 B2 GROUND PATTERN 1.08 0 0 .01n .01n 20n 011 R=-1
VFORCE__B3 B3 GROUND PATTERN 1.08 0 0 .01n .01n 20n 000 R=-1
VFORCE__A0 A0 GROUND PATTERN 1.08 0 0 .01n .01n 20n 111 R=-1
VFORCE__A1 A1 GROUND PATTERN 1.08 0 0 .01n .01n 20n 110 R=-1
VFORCE__A2 A2 GROUND PATTERN 1.08 0 0 .01n .01n 20n 101 R=-1
VFORCE__A3 A3 GROUND PATTERN 1.08 0 0 .01n .01n 20n 110 R=-1

* --- Global Outputs
.PROBE V SG

* --- Waveform Outputs
.PLOT DC V(COUT)
.PLOT TRAN V(COUT)

* --- Waveform Outputs for Group PROBES__S0
.PLOT DC V(S0) V(S1) V(S2) V(S3)
.PLOT TRAN V(S0) V(S1) V(S2) V(S3)

* --- Params
.TEMP 125

* --- Libsetup
.LIB KEY=MOS "$GENERIC13/models/lib.eldo" TT
.LIB KEY=MOS_33 "$GENERIC13/models/lib.eldo" TT_33
.LIB KEY=MOS_lvt "$GENERIC13/models/lib.eldo" TT_lvt
.LIB KEY=MOS_hvt "$GENERIC13/models/lib.eldo" TT_hvt
.LIB KEY=BIP "$GENERIC13/models/lib.eldo" TT_BIP
.LIB KEY=BIP_NPN "$GENERIC13/models/lib.eldo" TT_BIP_NPN
.LIB KEY=RES "$GENERIC13/models/lib.eldo" TT_RES
