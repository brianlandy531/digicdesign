.subckt PM_INV2_GROUND 1 2 16
-c0 22 0 0.15714f
-c1 19 0 0.281799f
-c2 13 0 0.329739f
-c3 10 0 0.228983f
-r4 17 19 0.327298
-r5 14 22 0.026824
-r6 14 16 0.100282
-r7 13 17 0.0453973
-r8 13 16 0.188169
-r9 8 22 0.0153724
-r10 8 10 0.29363
-r11 2 19 15.53
-r12 2 10 15.61
-r13 1 2 6.27522
.ends

.subckt PM_INV2_VOUT 1 3 8
-c0 18 0 0.537529f
-c1 16 0 0.10202f
-c2 13 0 0.09945f
-r5 8 11 0.0624
-r4 11 13 0.03584
-r3 16 18 0.0577135
-r6 5 13 0.0126293
-r7 5 18 1.16293
-r8 4 16 15.53
-r9 4 11 15.61
-r10 3 4 3.51923
-r11 1 4 6.01622
.ends

.subckt PM_INV2_VDD 1 3 12
-c0 21 0 0.16146f
-c1 15 0 0.103081f
-c2 9 0 0.251373f
-c3 8 0 0.23468f
-c4 7 0 0.0985f

-r5 13 15 0.0615211
-r6 10 21 0.0254635
-r7 10 12 0.044
-r8 9 13 0.0351279
-r9 9 12 0.173333
-r10 8 21 0.0168226
-r11 7 19 0.0611843
-r12 7 8 0.48186
-r13 1 3 3.44885
-r14 1 19 15.53
-r15 1 15 15.61
.ends

.subckt PM_INV2_VIN 4 8 12
-c0 12 0 0.1256f
-c1 10 0 0.166f
-c2 8 0 0.376634f
-c3 4 0 0.513364f

-r4 10 20 10.0225
-r5 10 18 9.82252
-r6 10 12 11.07
-r7 8 20 86.1538

-r8 4 18 133.077
.ends