* ELDO netlist generated with ICnet by 'bxl1703' on Thu Sep 12 2019 at 23:54:14

.CONNECT GROUND 0

*
* Globals.
*
.global GROUND

*
* MAIN CELL: Component pathname : $PYXIS_SPT/digicdesign/inv2
*
        M2 VOUT VIN GROUND N$50 nmos w=0.26u l=0.13u m=1 as=88.4f ad=88.4f
+  ps=0.94u pd=0.94u
        C1 VOUT GROUND 0
        M3 VOUT VIN VDD VDD pmos w=0.52u l=0.13u m=1 as=0.1768p ad=0.1768p
+  ps=1.2u pd=1.2u
*
.end
