* Example circuit file for simulating PEX

.OPTION DOTNODE
.HIER /

.INCLUDE "/home/bxl1703/Pyxis_SPT_HEP/ic_projects/Pyxis_SPT/digicdesign/4bitripplecarry/4bitripplecarry.cal/4bitripplecarry.pex.netlist"

.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_33
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_lwt
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_hwt
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_BIP
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_BIP_NPN
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo DIO
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo DIO_33
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo TT_RES
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/lib.eldo MOS_CAP
.LIB /home/bxl1703/Pyxis_SPT_HEP/ic_reflibs/tech_libs/generic13/models/res.spi res_t









* - Instantiate your parasitic netlist and add the load capacitor
** FORMAT : 
* XLAYOUT [all inputs as listed by the ".subckt" line in the included netlist, in the order that they appear there] [name of the subcircuit as listed in the included netlist]
XLAYOUT B0 CIN0 A0 S0 A1 B1 S1 B2 A2 S2 B3 A3 GROUND COUT S3 4BITRIPPLECARRY 

COUT S0 0 120f
COUT S1 0 120f
COUT S2 0 120f
COUT S3 0 120f
COUT COUT 0 120f

* - Analysis Setup - DC sweep
* FORMAT : .DC [name] [low] [high] [step]
* .DC VFORCE__VIN 0 1.08 0.01

* - Analysis Setup - Trans
* FORMAT : .TRAN [start time] [end time] [time step]
.TRAN 0 10000n 0.001n

* --- Forces
* FORMAT -- PULSE : [name] [port] [reference (0 means ground)] PULSE [low] [high] [delay] [fall time] [rise time] [pulse width] [period]
*
* FORMAT -- DC    : [name] [port] [reference (0 means ground)] DC [voltage]
*
** VFORCE__Vin VIN 0 PULSE (0 1.08 100n 0.1n 0.1n 50n 200n)

VFORCE__VDD VDD 0 DC 1.08
VFORCE__GROUND GROUND 0 DC 0

VFORCE__B0 B0 0 pattern 1.08 0 50n .01n .01n 100n 011 R
VFORCE__B1 B1 0 pattern 1.08 0 50n .01n .01n 100n 010 R
VFORCE__B2 B2 0 pattern 1.08 0 50n .01n .01n 100n 011 R
VFORCE__B3 B3 0 pattern 1.08 0 50n .01n .01n 100n 000 R


VFORCE__A0 A0 0 pattern 1.08 0 50n .01n .01n 100n 111 R
VFORCE__A1 A1 0 pattern 1.08 0 50n .01n .01n 100n 110 R
VFORCE__A2 A2 0 pattern 1.08 0 50n .01n .01n 100n 101 R
VFORCE__A3 A3 0 pattern 1.08 0 50n .01n .01n 100n 110 R


VFORCE__CIN0 CIN0 0 pattern 1.08 0 50n .01n .01n 100n 101 R

* --- Waveform Outputs
*.PLOT DC V(VIN)
*.PLOT DC V(VOUT)
.PLOT TRAN V(CIN0)


.PLOT TRAN V(COUT)

.PLOT TRAN V(A0)
.PLOT TRAN V(A1)
.PLOT TRAN V(A2)
.PLOT TRAN V(A3)

.PLOT TRAN V(B0)
.PLOT TRAN V(B1)
.PLOT TRAN V(B2)
.PLOT TRAN V(B3)

.PLOT TRAN V(S0)
.PLOT TRAN V(S1)
.PLOT TRAN V(S2)
.PLOT TRAN V(S3)



* --- Params
.TEMP 125


